# This file is SVn file which
# is having evn variable

Cloude=azure
Resource=ec2
Name=Test
enveronment=Test


Cloude=azure
Resource=ec2
Name=Test
enveronment=Test



